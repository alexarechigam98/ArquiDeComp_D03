
//1.Definicion del modulo y sus I/O
//Dentro del parentesis se define los I/O
module _and(input a, input b, output c);
//2.Definen cables o componenetes internos
//NA
//3. Asignaciones, instancias, conexiones

assign c = a & b;

endmodule